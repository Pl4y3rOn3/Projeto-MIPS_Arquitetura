// Verilog code for instruction memory
 module instr_mem          // a synthesisable rom implementation  
 (  
      input [31:0] pc, //Address PC 
      output wire [31:0] instruction //i_out
 );  
      wire [4 : 0] rom_addr = pc[5 : 1];  //Index
		
      reg [31:0] rom [31:0];  //32 intruções de 32 bits
      initial  
      begin  
                rom[0] = 32'b00000000000000000000000000000000; //
                rom[1] = 32'b00000000000000000000000000000000; //
                rom[2] = 32'b00000000000000000000000000000000; //
                rom[3] = 32'b00000000000000000000000000000000; //
                rom[4] = 32'b00000000000000000000000000000000; //
                rom[5] = 32'b00000000000000000000000000000000; //
					 rom[6] = 32'b00000000000000000000000000000000; //
                rom[7] = 32'b00000000000000000000000000000000; //
                rom[8] = 32'b00000000000000000000000000000000; //
                rom[9] = 32'b00000000000000000000000000000000; //
                rom[10] = 32'b00000000000000000000000000000000;// 
                rom[11] = 32'b00000000000000000000000000000000;//
					 rom[12] = 32'b00000000000000000000000000000000;//
                rom[13] = 32'b00000000000000000000000000000000;//
                rom[14] = 32'b00000000000000000000000000000000;//
                rom[15] = 32'b00000000000000000000000000000000;//
                rom[16] = 32'b00000000000000000000000000000000;//
                rom[17] = 32'b00000000000000000000000000000000;//
					 rom[18] = 32'b00000000000000000000000000000000;//	
                rom[19] = 32'b00000000000000000000000000000000;//
                rom[20] = 32'b00000000000000000000000000000000;//
                rom[21] = 32'b00000000000000000000000000000000;//
                rom[22] = 32'b00000000000000000000000000000000;//
                rom[23] = 32'b00000000000000000000000000000000;//
					 rom[24] = 32'b00000000000000000000000000000000;//	
                rom[25] = 32'b00000000000000000000000000000000;//  
                rom[26] = 32'b00000000000000000000000000000000;//
                rom[27] = 32'b00000000000000000000000000000000;  
                rom[28] = 32'b00000000000000000000000000000000;  
                rom[29] = 32'b00000000000000000000000000000000;
					 rom[30] = 32'b00000000000000000000000000000000;  	
                rom[31] = 32'b00000000000000000000000000000000;  
                  
      end  
      assign instruction = (pc[31:0] < 64 )? rom[rom_addr[4:0]]: 32'd0;  
 endmodule 